Patrol|Address1|Address2|Address3|Address4|Address5|
09|ASIAN CENTRE, 50|ABBEY ROAD||||
